
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'haedd12c0;
    ram_cell[       1] = 32'h0;  // 32'hd7342c94;
    ram_cell[       2] = 32'h0;  // 32'h545494db;
    ram_cell[       3] = 32'h0;  // 32'h669f25fe;
    ram_cell[       4] = 32'h0;  // 32'h78f6b773;
    ram_cell[       5] = 32'h0;  // 32'heb20963d;
    ram_cell[       6] = 32'h0;  // 32'h8be5a4dd;
    ram_cell[       7] = 32'h0;  // 32'h5411bd21;
    ram_cell[       8] = 32'h0;  // 32'habdfabea;
    ram_cell[       9] = 32'h0;  // 32'hfa8770c3;
    ram_cell[      10] = 32'h0;  // 32'h7777a3df;
    ram_cell[      11] = 32'h0;  // 32'hf010a849;
    ram_cell[      12] = 32'h0;  // 32'h0652408f;
    ram_cell[      13] = 32'h0;  // 32'h011c5306;
    ram_cell[      14] = 32'h0;  // 32'h0d6f75ba;
    ram_cell[      15] = 32'h0;  // 32'h392d86e9;
    ram_cell[      16] = 32'h0;  // 32'h6da2629d;
    ram_cell[      17] = 32'h0;  // 32'h1093284b;
    ram_cell[      18] = 32'h0;  // 32'h5454bdac;
    ram_cell[      19] = 32'h0;  // 32'hefc8dde6;
    ram_cell[      20] = 32'h0;  // 32'he0b82137;
    ram_cell[      21] = 32'h0;  // 32'h1c6a2e70;
    ram_cell[      22] = 32'h0;  // 32'h66b79e0e;
    ram_cell[      23] = 32'h0;  // 32'hb8ad8290;
    ram_cell[      24] = 32'h0;  // 32'h8af5c372;
    ram_cell[      25] = 32'h0;  // 32'he014de60;
    ram_cell[      26] = 32'h0;  // 32'hf6456adf;
    ram_cell[      27] = 32'h0;  // 32'h65cde318;
    ram_cell[      28] = 32'h0;  // 32'hf178ebd9;
    ram_cell[      29] = 32'h0;  // 32'had9205a5;
    ram_cell[      30] = 32'h0;  // 32'hf11a1991;
    ram_cell[      31] = 32'h0;  // 32'hb3c45e2b;
    ram_cell[      32] = 32'h0;  // 32'h9c8b0a9c;
    ram_cell[      33] = 32'h0;  // 32'h52506420;
    ram_cell[      34] = 32'h0;  // 32'h71fd6f29;
    ram_cell[      35] = 32'h0;  // 32'h570f8765;
    ram_cell[      36] = 32'h0;  // 32'hdde0bb16;
    ram_cell[      37] = 32'h0;  // 32'hdfc536e9;
    ram_cell[      38] = 32'h0;  // 32'h926300e7;
    ram_cell[      39] = 32'h0;  // 32'he853c002;
    ram_cell[      40] = 32'h0;  // 32'hd97271b8;
    ram_cell[      41] = 32'h0;  // 32'h180c75cb;
    ram_cell[      42] = 32'h0;  // 32'hcae8cb6e;
    ram_cell[      43] = 32'h0;  // 32'he8933d46;
    ram_cell[      44] = 32'h0;  // 32'hdfb87915;
    ram_cell[      45] = 32'h0;  // 32'ha1e729c0;
    ram_cell[      46] = 32'h0;  // 32'h32077f12;
    ram_cell[      47] = 32'h0;  // 32'ha2f56b86;
    ram_cell[      48] = 32'h0;  // 32'he37eaad5;
    ram_cell[      49] = 32'h0;  // 32'h48e7a14a;
    ram_cell[      50] = 32'h0;  // 32'hf4de76de;
    ram_cell[      51] = 32'h0;  // 32'heed69ffd;
    ram_cell[      52] = 32'h0;  // 32'h1b413933;
    ram_cell[      53] = 32'h0;  // 32'h8cacf01c;
    ram_cell[      54] = 32'h0;  // 32'h07cb553d;
    ram_cell[      55] = 32'h0;  // 32'hec4cd526;
    ram_cell[      56] = 32'h0;  // 32'h5246daaa;
    ram_cell[      57] = 32'h0;  // 32'h100274de;
    ram_cell[      58] = 32'h0;  // 32'h6418a981;
    ram_cell[      59] = 32'h0;  // 32'h9423f426;
    ram_cell[      60] = 32'h0;  // 32'h191751b0;
    ram_cell[      61] = 32'h0;  // 32'hce4bf658;
    ram_cell[      62] = 32'h0;  // 32'hf87ed7c3;
    ram_cell[      63] = 32'h0;  // 32'h9d239cde;
    ram_cell[      64] = 32'h0;  // 32'h8a6a2deb;
    ram_cell[      65] = 32'h0;  // 32'h0c0fc23e;
    ram_cell[      66] = 32'h0;  // 32'h21059f66;
    ram_cell[      67] = 32'h0;  // 32'h836738c4;
    ram_cell[      68] = 32'h0;  // 32'h35f96165;
    ram_cell[      69] = 32'h0;  // 32'h6e124411;
    ram_cell[      70] = 32'h0;  // 32'h2bf91aaa;
    ram_cell[      71] = 32'h0;  // 32'hcf4f9499;
    ram_cell[      72] = 32'h0;  // 32'h4fadeaaf;
    ram_cell[      73] = 32'h0;  // 32'h544d9029;
    ram_cell[      74] = 32'h0;  // 32'h597f12b9;
    ram_cell[      75] = 32'h0;  // 32'h24d5ee50;
    ram_cell[      76] = 32'h0;  // 32'h9b287306;
    ram_cell[      77] = 32'h0;  // 32'h6b853495;
    ram_cell[      78] = 32'h0;  // 32'h82eedc64;
    ram_cell[      79] = 32'h0;  // 32'hd8bade8a;
    ram_cell[      80] = 32'h0;  // 32'h7eebba18;
    ram_cell[      81] = 32'h0;  // 32'h45999c53;
    ram_cell[      82] = 32'h0;  // 32'ha98557ca;
    ram_cell[      83] = 32'h0;  // 32'h94efeab1;
    ram_cell[      84] = 32'h0;  // 32'hefcd1ebb;
    ram_cell[      85] = 32'h0;  // 32'h1b98c312;
    ram_cell[      86] = 32'h0;  // 32'haa29edd1;
    ram_cell[      87] = 32'h0;  // 32'h4d84ae04;
    ram_cell[      88] = 32'h0;  // 32'hdbb435e4;
    ram_cell[      89] = 32'h0;  // 32'h87d541a6;
    ram_cell[      90] = 32'h0;  // 32'ha3e4a34d;
    ram_cell[      91] = 32'h0;  // 32'h3f504b92;
    ram_cell[      92] = 32'h0;  // 32'h9d80394a;
    ram_cell[      93] = 32'h0;  // 32'h6208fef8;
    ram_cell[      94] = 32'h0;  // 32'hacf0cfb3;
    ram_cell[      95] = 32'h0;  // 32'hb43fcda0;
    ram_cell[      96] = 32'h0;  // 32'hd1963aba;
    ram_cell[      97] = 32'h0;  // 32'had1439b3;
    ram_cell[      98] = 32'h0;  // 32'h4234c1a5;
    ram_cell[      99] = 32'h0;  // 32'h6228d79f;
    ram_cell[     100] = 32'h0;  // 32'h459c9592;
    ram_cell[     101] = 32'h0;  // 32'h39a261ef;
    ram_cell[     102] = 32'h0;  // 32'hdd7b7bbf;
    ram_cell[     103] = 32'h0;  // 32'h2d2e3ef9;
    ram_cell[     104] = 32'h0;  // 32'h82dd1dc1;
    ram_cell[     105] = 32'h0;  // 32'h90ca9664;
    ram_cell[     106] = 32'h0;  // 32'h4dc77fe6;
    ram_cell[     107] = 32'h0;  // 32'h6da55b9c;
    ram_cell[     108] = 32'h0;  // 32'hb1448a31;
    ram_cell[     109] = 32'h0;  // 32'h18be7598;
    ram_cell[     110] = 32'h0;  // 32'h6d15524e;
    ram_cell[     111] = 32'h0;  // 32'h1fcb5936;
    ram_cell[     112] = 32'h0;  // 32'hc2b6288d;
    ram_cell[     113] = 32'h0;  // 32'h7c72aa40;
    ram_cell[     114] = 32'h0;  // 32'h6893b995;
    ram_cell[     115] = 32'h0;  // 32'h09ffb959;
    ram_cell[     116] = 32'h0;  // 32'h615e4c93;
    ram_cell[     117] = 32'h0;  // 32'hbdc03e75;
    ram_cell[     118] = 32'h0;  // 32'h99c39a38;
    ram_cell[     119] = 32'h0;  // 32'hf6d7cfb7;
    ram_cell[     120] = 32'h0;  // 32'hc3575b1c;
    ram_cell[     121] = 32'h0;  // 32'hef1f2c05;
    ram_cell[     122] = 32'h0;  // 32'h6e28eb69;
    ram_cell[     123] = 32'h0;  // 32'h1b43aa38;
    ram_cell[     124] = 32'h0;  // 32'h5042461b;
    ram_cell[     125] = 32'h0;  // 32'h53acce8a;
    ram_cell[     126] = 32'h0;  // 32'he20a616c;
    ram_cell[     127] = 32'h0;  // 32'h5abfcebf;
    ram_cell[     128] = 32'h0;  // 32'h8c4768c8;
    ram_cell[     129] = 32'h0;  // 32'hb6981c99;
    ram_cell[     130] = 32'h0;  // 32'hacefd645;
    ram_cell[     131] = 32'h0;  // 32'h27f7d9be;
    ram_cell[     132] = 32'h0;  // 32'hbf73a2f6;
    ram_cell[     133] = 32'h0;  // 32'hf16d4bc9;
    ram_cell[     134] = 32'h0;  // 32'h01270019;
    ram_cell[     135] = 32'h0;  // 32'h66b5f008;
    ram_cell[     136] = 32'h0;  // 32'h56d81f43;
    ram_cell[     137] = 32'h0;  // 32'h2f9e4d73;
    ram_cell[     138] = 32'h0;  // 32'h3aadbf69;
    ram_cell[     139] = 32'h0;  // 32'h392a8c40;
    ram_cell[     140] = 32'h0;  // 32'h8d5fd25e;
    ram_cell[     141] = 32'h0;  // 32'h50f75ad6;
    ram_cell[     142] = 32'h0;  // 32'h7328aaef;
    ram_cell[     143] = 32'h0;  // 32'h30f4ba4e;
    ram_cell[     144] = 32'h0;  // 32'ha43f702a;
    ram_cell[     145] = 32'h0;  // 32'h90d4f31c;
    ram_cell[     146] = 32'h0;  // 32'h64432db7;
    ram_cell[     147] = 32'h0;  // 32'h5951ebb8;
    ram_cell[     148] = 32'h0;  // 32'hce22c5a5;
    ram_cell[     149] = 32'h0;  // 32'hafa7bc13;
    ram_cell[     150] = 32'h0;  // 32'hc77727a5;
    ram_cell[     151] = 32'h0;  // 32'h27fb05f2;
    ram_cell[     152] = 32'h0;  // 32'ha9de99bb;
    ram_cell[     153] = 32'h0;  // 32'h993d8a2e;
    ram_cell[     154] = 32'h0;  // 32'hc27b5ae3;
    ram_cell[     155] = 32'h0;  // 32'hd98c6a6f;
    ram_cell[     156] = 32'h0;  // 32'h16c345e9;
    ram_cell[     157] = 32'h0;  // 32'hd28819d4;
    ram_cell[     158] = 32'h0;  // 32'h73af92a5;
    ram_cell[     159] = 32'h0;  // 32'h0ea1c750;
    ram_cell[     160] = 32'h0;  // 32'hd7f9fac3;
    ram_cell[     161] = 32'h0;  // 32'h1f6a0ac1;
    ram_cell[     162] = 32'h0;  // 32'haf4cfd38;
    ram_cell[     163] = 32'h0;  // 32'hff9d4329;
    ram_cell[     164] = 32'h0;  // 32'h0c784a42;
    ram_cell[     165] = 32'h0;  // 32'h01260c6e;
    ram_cell[     166] = 32'h0;  // 32'h4b74f56e;
    ram_cell[     167] = 32'h0;  // 32'h841935a8;
    ram_cell[     168] = 32'h0;  // 32'hefc829ec;
    ram_cell[     169] = 32'h0;  // 32'h895dab17;
    ram_cell[     170] = 32'h0;  // 32'h2036d238;
    ram_cell[     171] = 32'h0;  // 32'h4bfdaf12;
    ram_cell[     172] = 32'h0;  // 32'h188a9844;
    ram_cell[     173] = 32'h0;  // 32'h7792efba;
    ram_cell[     174] = 32'h0;  // 32'h5d35c1ed;
    ram_cell[     175] = 32'h0;  // 32'h012ef917;
    ram_cell[     176] = 32'h0;  // 32'h80ee7ee3;
    ram_cell[     177] = 32'h0;  // 32'ha611a9f2;
    ram_cell[     178] = 32'h0;  // 32'heafac231;
    ram_cell[     179] = 32'h0;  // 32'h1726e9bb;
    ram_cell[     180] = 32'h0;  // 32'h8d457e77;
    ram_cell[     181] = 32'h0;  // 32'h17dda4f7;
    ram_cell[     182] = 32'h0;  // 32'h72903b04;
    ram_cell[     183] = 32'h0;  // 32'ha4ec0432;
    ram_cell[     184] = 32'h0;  // 32'h029d3e11;
    ram_cell[     185] = 32'h0;  // 32'h34077bcf;
    ram_cell[     186] = 32'h0;  // 32'h290e82b7;
    ram_cell[     187] = 32'h0;  // 32'h8d5f459d;
    ram_cell[     188] = 32'h0;  // 32'h11074363;
    ram_cell[     189] = 32'h0;  // 32'h908fc848;
    ram_cell[     190] = 32'h0;  // 32'h75069133;
    ram_cell[     191] = 32'h0;  // 32'h0547115d;
    ram_cell[     192] = 32'h0;  // 32'h5cdcff5f;
    ram_cell[     193] = 32'h0;  // 32'hdf9058cd;
    ram_cell[     194] = 32'h0;  // 32'h0154eb5f;
    ram_cell[     195] = 32'h0;  // 32'h8bea56db;
    ram_cell[     196] = 32'h0;  // 32'h03be5c0c;
    ram_cell[     197] = 32'h0;  // 32'hc88ada8e;
    ram_cell[     198] = 32'h0;  // 32'hbafb32c9;
    ram_cell[     199] = 32'h0;  // 32'h1a5ef4f9;
    ram_cell[     200] = 32'h0;  // 32'h25c94c82;
    ram_cell[     201] = 32'h0;  // 32'h2ba2ecbd;
    ram_cell[     202] = 32'h0;  // 32'h74ace757;
    ram_cell[     203] = 32'h0;  // 32'hb5b9a700;
    ram_cell[     204] = 32'h0;  // 32'hc759ee59;
    ram_cell[     205] = 32'h0;  // 32'hdd88b757;
    ram_cell[     206] = 32'h0;  // 32'h659dbf35;
    ram_cell[     207] = 32'h0;  // 32'hb884b237;
    ram_cell[     208] = 32'h0;  // 32'h652805d1;
    ram_cell[     209] = 32'h0;  // 32'h40beaf12;
    ram_cell[     210] = 32'h0;  // 32'h0005eedc;
    ram_cell[     211] = 32'h0;  // 32'h667156d1;
    ram_cell[     212] = 32'h0;  // 32'hc4b240cb;
    ram_cell[     213] = 32'h0;  // 32'h6a56f1a8;
    ram_cell[     214] = 32'h0;  // 32'h90f40761;
    ram_cell[     215] = 32'h0;  // 32'h1373658d;
    ram_cell[     216] = 32'h0;  // 32'h4482b4d5;
    ram_cell[     217] = 32'h0;  // 32'ha09140bd;
    ram_cell[     218] = 32'h0;  // 32'h8d60a107;
    ram_cell[     219] = 32'h0;  // 32'h34e8622f;
    ram_cell[     220] = 32'h0;  // 32'h791d2e52;
    ram_cell[     221] = 32'h0;  // 32'h0feb9468;
    ram_cell[     222] = 32'h0;  // 32'h0131c92a;
    ram_cell[     223] = 32'h0;  // 32'hff39d865;
    ram_cell[     224] = 32'h0;  // 32'h35892c36;
    ram_cell[     225] = 32'h0;  // 32'h3d76b0c6;
    ram_cell[     226] = 32'h0;  // 32'h920c0d43;
    ram_cell[     227] = 32'h0;  // 32'he5ee94d0;
    ram_cell[     228] = 32'h0;  // 32'hb926ce1f;
    ram_cell[     229] = 32'h0;  // 32'h033e4cf6;
    ram_cell[     230] = 32'h0;  // 32'h8e433ba7;
    ram_cell[     231] = 32'h0;  // 32'h90ffec4f;
    ram_cell[     232] = 32'h0;  // 32'h3843228c;
    ram_cell[     233] = 32'h0;  // 32'hf4ca03da;
    ram_cell[     234] = 32'h0;  // 32'h70c4bae5;
    ram_cell[     235] = 32'h0;  // 32'h96d1461e;
    ram_cell[     236] = 32'h0;  // 32'h72b91de4;
    ram_cell[     237] = 32'h0;  // 32'ha1d824b3;
    ram_cell[     238] = 32'h0;  // 32'hdfc0f6db;
    ram_cell[     239] = 32'h0;  // 32'h494082dd;
    ram_cell[     240] = 32'h0;  // 32'h26ee1d1d;
    ram_cell[     241] = 32'h0;  // 32'h77e3c4e0;
    ram_cell[     242] = 32'h0;  // 32'h21c3a759;
    ram_cell[     243] = 32'h0;  // 32'h2afc95b0;
    ram_cell[     244] = 32'h0;  // 32'h3fd348d6;
    ram_cell[     245] = 32'h0;  // 32'h595a2254;
    ram_cell[     246] = 32'h0;  // 32'h57c66fc0;
    ram_cell[     247] = 32'h0;  // 32'heb420f61;
    ram_cell[     248] = 32'h0;  // 32'h24df786f;
    ram_cell[     249] = 32'h0;  // 32'h6ca63250;
    ram_cell[     250] = 32'h0;  // 32'h65200d0a;
    ram_cell[     251] = 32'h0;  // 32'he8ca8497;
    ram_cell[     252] = 32'h0;  // 32'h315c0d90;
    ram_cell[     253] = 32'h0;  // 32'h998895b1;
    ram_cell[     254] = 32'h0;  // 32'hc212dbc6;
    ram_cell[     255] = 32'h0;  // 32'hc21dcc2e;
    // src matrix A
    ram_cell[     256] = 32'hcb27a532;
    ram_cell[     257] = 32'hbf2d0df6;
    ram_cell[     258] = 32'hdf680697;
    ram_cell[     259] = 32'h430dc3c6;
    ram_cell[     260] = 32'h3c560a86;
    ram_cell[     261] = 32'h659f7215;
    ram_cell[     262] = 32'h092b27f3;
    ram_cell[     263] = 32'h69e72c6a;
    ram_cell[     264] = 32'h853a5c1a;
    ram_cell[     265] = 32'h5aa864c6;
    ram_cell[     266] = 32'h795dc057;
    ram_cell[     267] = 32'h91c195f5;
    ram_cell[     268] = 32'h10a058ed;
    ram_cell[     269] = 32'h10bed988;
    ram_cell[     270] = 32'hb2ea7690;
    ram_cell[     271] = 32'hc9dbdef6;
    ram_cell[     272] = 32'h20f8ec6d;
    ram_cell[     273] = 32'h94b66711;
    ram_cell[     274] = 32'hba7dc859;
    ram_cell[     275] = 32'hb55768bc;
    ram_cell[     276] = 32'hc4475ff6;
    ram_cell[     277] = 32'h9bad9449;
    ram_cell[     278] = 32'h93650ac6;
    ram_cell[     279] = 32'h85f8eb49;
    ram_cell[     280] = 32'he938ca90;
    ram_cell[     281] = 32'h3f25b606;
    ram_cell[     282] = 32'h52774413;
    ram_cell[     283] = 32'h388da401;
    ram_cell[     284] = 32'h76881e0e;
    ram_cell[     285] = 32'hb163e811;
    ram_cell[     286] = 32'hbd49cbd1;
    ram_cell[     287] = 32'h84c52b65;
    ram_cell[     288] = 32'h133e46dd;
    ram_cell[     289] = 32'h09d55412;
    ram_cell[     290] = 32'h71425567;
    ram_cell[     291] = 32'ha25d40e0;
    ram_cell[     292] = 32'h1b8d1a29;
    ram_cell[     293] = 32'h8e1c4b82;
    ram_cell[     294] = 32'h8ac05927;
    ram_cell[     295] = 32'h4369a56d;
    ram_cell[     296] = 32'hc2364888;
    ram_cell[     297] = 32'hdcf953ee;
    ram_cell[     298] = 32'h165ea9a0;
    ram_cell[     299] = 32'ha4b3cc8f;
    ram_cell[     300] = 32'hd2aa268c;
    ram_cell[     301] = 32'hb3a45811;
    ram_cell[     302] = 32'hbbe90e14;
    ram_cell[     303] = 32'hbc14a335;
    ram_cell[     304] = 32'h8195d061;
    ram_cell[     305] = 32'h78b59299;
    ram_cell[     306] = 32'h80f28618;
    ram_cell[     307] = 32'h2fa068ae;
    ram_cell[     308] = 32'hb77c9cec;
    ram_cell[     309] = 32'h943f308e;
    ram_cell[     310] = 32'h6427e856;
    ram_cell[     311] = 32'heaf114ee;
    ram_cell[     312] = 32'h8e7d8ecc;
    ram_cell[     313] = 32'h23b94d55;
    ram_cell[     314] = 32'h015bae34;
    ram_cell[     315] = 32'h27f2f290;
    ram_cell[     316] = 32'hc6ede56f;
    ram_cell[     317] = 32'hb5b015e5;
    ram_cell[     318] = 32'hf3e4ede3;
    ram_cell[     319] = 32'h96d2a175;
    ram_cell[     320] = 32'ha176b87d;
    ram_cell[     321] = 32'hf3c53546;
    ram_cell[     322] = 32'h26500d86;
    ram_cell[     323] = 32'h8e41d26b;
    ram_cell[     324] = 32'h33129620;
    ram_cell[     325] = 32'h1231b865;
    ram_cell[     326] = 32'ha72bfc34;
    ram_cell[     327] = 32'h9ee529a0;
    ram_cell[     328] = 32'h185e6ac3;
    ram_cell[     329] = 32'h4e6a2bae;
    ram_cell[     330] = 32'h08a53659;
    ram_cell[     331] = 32'h280c82db;
    ram_cell[     332] = 32'h5cad5948;
    ram_cell[     333] = 32'hb8fc67e3;
    ram_cell[     334] = 32'h19d7b2fe;
    ram_cell[     335] = 32'hfc33f3b1;
    ram_cell[     336] = 32'h72069ca9;
    ram_cell[     337] = 32'hb0731d44;
    ram_cell[     338] = 32'ha79632d2;
    ram_cell[     339] = 32'h1a442ddf;
    ram_cell[     340] = 32'h13af3d6c;
    ram_cell[     341] = 32'h0d558d3c;
    ram_cell[     342] = 32'h831d0f0b;
    ram_cell[     343] = 32'h5297ef89;
    ram_cell[     344] = 32'hf568d433;
    ram_cell[     345] = 32'h6cd9d6b4;
    ram_cell[     346] = 32'h7626e1d1;
    ram_cell[     347] = 32'h9e88d94d;
    ram_cell[     348] = 32'h3ab3523d;
    ram_cell[     349] = 32'h206247df;
    ram_cell[     350] = 32'h33675be0;
    ram_cell[     351] = 32'h14a6a544;
    ram_cell[     352] = 32'he76ce7eb;
    ram_cell[     353] = 32'hd34c2527;
    ram_cell[     354] = 32'h694b34f9;
    ram_cell[     355] = 32'hc428566f;
    ram_cell[     356] = 32'h7f53cd86;
    ram_cell[     357] = 32'ha1318781;
    ram_cell[     358] = 32'h0a028530;
    ram_cell[     359] = 32'h9d9940a7;
    ram_cell[     360] = 32'hee5f6edc;
    ram_cell[     361] = 32'h116556b8;
    ram_cell[     362] = 32'hf01056b1;
    ram_cell[     363] = 32'hecd35ebf;
    ram_cell[     364] = 32'h2afa5e9e;
    ram_cell[     365] = 32'h7512055a;
    ram_cell[     366] = 32'hc4804340;
    ram_cell[     367] = 32'h5000f03d;
    ram_cell[     368] = 32'hf2510fe4;
    ram_cell[     369] = 32'h3e896391;
    ram_cell[     370] = 32'hee5091b4;
    ram_cell[     371] = 32'hfe4d30ff;
    ram_cell[     372] = 32'h370fc498;
    ram_cell[     373] = 32'h5236a931;
    ram_cell[     374] = 32'h84035092;
    ram_cell[     375] = 32'h47238ec9;
    ram_cell[     376] = 32'he5b28199;
    ram_cell[     377] = 32'h01453186;
    ram_cell[     378] = 32'hd4968678;
    ram_cell[     379] = 32'hacb2d440;
    ram_cell[     380] = 32'hdfe78ef6;
    ram_cell[     381] = 32'h9fda525a;
    ram_cell[     382] = 32'h367cc8f2;
    ram_cell[     383] = 32'h561dba1c;
    ram_cell[     384] = 32'h6a62252e;
    ram_cell[     385] = 32'h45b0edc2;
    ram_cell[     386] = 32'hba34655c;
    ram_cell[     387] = 32'h782c0ab0;
    ram_cell[     388] = 32'h9b4d43b9;
    ram_cell[     389] = 32'h421217d1;
    ram_cell[     390] = 32'h0bb5cce5;
    ram_cell[     391] = 32'h2952a60a;
    ram_cell[     392] = 32'h2eed8a6c;
    ram_cell[     393] = 32'h9eaf2943;
    ram_cell[     394] = 32'hf1eb79ab;
    ram_cell[     395] = 32'he5ec431a;
    ram_cell[     396] = 32'h23b85a30;
    ram_cell[     397] = 32'h5483901a;
    ram_cell[     398] = 32'hea5e2725;
    ram_cell[     399] = 32'h6d356513;
    ram_cell[     400] = 32'he91a6375;
    ram_cell[     401] = 32'h2d43f4be;
    ram_cell[     402] = 32'he098a666;
    ram_cell[     403] = 32'h1db69ddf;
    ram_cell[     404] = 32'hea2eeecb;
    ram_cell[     405] = 32'h9a64de12;
    ram_cell[     406] = 32'h03376ec3;
    ram_cell[     407] = 32'h75f4653b;
    ram_cell[     408] = 32'h9ca0b205;
    ram_cell[     409] = 32'h10459933;
    ram_cell[     410] = 32'hb7852518;
    ram_cell[     411] = 32'hd9688bea;
    ram_cell[     412] = 32'h02f1d1ad;
    ram_cell[     413] = 32'hdfb74866;
    ram_cell[     414] = 32'hf1ed853b;
    ram_cell[     415] = 32'hb14a066b;
    ram_cell[     416] = 32'h5e3e6193;
    ram_cell[     417] = 32'h5be34017;
    ram_cell[     418] = 32'hb508c4a5;
    ram_cell[     419] = 32'h4b3bcdc4;
    ram_cell[     420] = 32'h61249b7e;
    ram_cell[     421] = 32'h22f88fc3;
    ram_cell[     422] = 32'hab362ec2;
    ram_cell[     423] = 32'h4e8d592c;
    ram_cell[     424] = 32'h8de673b5;
    ram_cell[     425] = 32'h417c62da;
    ram_cell[     426] = 32'hf2c805da;
    ram_cell[     427] = 32'h4284ec6e;
    ram_cell[     428] = 32'hf038a56f;
    ram_cell[     429] = 32'hcfcac79b;
    ram_cell[     430] = 32'hef58d0fd;
    ram_cell[     431] = 32'h6fa6c695;
    ram_cell[     432] = 32'hf1610849;
    ram_cell[     433] = 32'h444153a3;
    ram_cell[     434] = 32'h433e726b;
    ram_cell[     435] = 32'h2fc4fc7d;
    ram_cell[     436] = 32'h2e4300c0;
    ram_cell[     437] = 32'hf6d7ddf6;
    ram_cell[     438] = 32'he6416f82;
    ram_cell[     439] = 32'h50a92b73;
    ram_cell[     440] = 32'he445d4a5;
    ram_cell[     441] = 32'h539326b1;
    ram_cell[     442] = 32'hd89972d8;
    ram_cell[     443] = 32'h4b36d777;
    ram_cell[     444] = 32'hc54e6d5c;
    ram_cell[     445] = 32'hdec765ec;
    ram_cell[     446] = 32'h656c5cae;
    ram_cell[     447] = 32'he0811d2a;
    ram_cell[     448] = 32'h838a4d40;
    ram_cell[     449] = 32'h3bcd4d61;
    ram_cell[     450] = 32'h85cecfe2;
    ram_cell[     451] = 32'hf48cda8b;
    ram_cell[     452] = 32'hd1a2a92a;
    ram_cell[     453] = 32'hb4eca359;
    ram_cell[     454] = 32'h01c08ec7;
    ram_cell[     455] = 32'h99422435;
    ram_cell[     456] = 32'h0db8689b;
    ram_cell[     457] = 32'h5a378eba;
    ram_cell[     458] = 32'h19cbee41;
    ram_cell[     459] = 32'hdcc8f4d9;
    ram_cell[     460] = 32'he247456e;
    ram_cell[     461] = 32'hf4996326;
    ram_cell[     462] = 32'h8fad1a0a;
    ram_cell[     463] = 32'h3a7efd7f;
    ram_cell[     464] = 32'heb1ffe81;
    ram_cell[     465] = 32'hf8919019;
    ram_cell[     466] = 32'h852586d5;
    ram_cell[     467] = 32'hc5e6efb5;
    ram_cell[     468] = 32'h737726cb;
    ram_cell[     469] = 32'h73b989de;
    ram_cell[     470] = 32'h185ba38e;
    ram_cell[     471] = 32'hdb454ff2;
    ram_cell[     472] = 32'h36a4cf50;
    ram_cell[     473] = 32'hcb73666c;
    ram_cell[     474] = 32'h2b36e262;
    ram_cell[     475] = 32'h37ff77b9;
    ram_cell[     476] = 32'h7619359f;
    ram_cell[     477] = 32'h1a659eca;
    ram_cell[     478] = 32'h9eddaa84;
    ram_cell[     479] = 32'hc63e30d4;
    ram_cell[     480] = 32'hb3632fa8;
    ram_cell[     481] = 32'h88c4eb96;
    ram_cell[     482] = 32'hd293729e;
    ram_cell[     483] = 32'h08daa593;
    ram_cell[     484] = 32'hb96c9a8d;
    ram_cell[     485] = 32'h8813c185;
    ram_cell[     486] = 32'hecf282bb;
    ram_cell[     487] = 32'h43beb6af;
    ram_cell[     488] = 32'hf09ca535;
    ram_cell[     489] = 32'h2d645433;
    ram_cell[     490] = 32'h3088479c;
    ram_cell[     491] = 32'h429159ca;
    ram_cell[     492] = 32'haedd173d;
    ram_cell[     493] = 32'hddc8d856;
    ram_cell[     494] = 32'hba770adb;
    ram_cell[     495] = 32'hea9d567b;
    ram_cell[     496] = 32'h95c9843d;
    ram_cell[     497] = 32'hf33c1aef;
    ram_cell[     498] = 32'h0b098cf1;
    ram_cell[     499] = 32'h89ddb398;
    ram_cell[     500] = 32'h2c738d63;
    ram_cell[     501] = 32'h2d724202;
    ram_cell[     502] = 32'hb040cd13;
    ram_cell[     503] = 32'hac5d4050;
    ram_cell[     504] = 32'had44bce8;
    ram_cell[     505] = 32'h930458c6;
    ram_cell[     506] = 32'ha0c9aad2;
    ram_cell[     507] = 32'ha5474319;
    ram_cell[     508] = 32'h28979708;
    ram_cell[     509] = 32'h3bd603ba;
    ram_cell[     510] = 32'h2d7e5944;
    ram_cell[     511] = 32'h1b3ec3f6;
    // src matrix B
    ram_cell[     512] = 32'h8f854653;
    ram_cell[     513] = 32'h878ba0be;
    ram_cell[     514] = 32'h6075afe3;
    ram_cell[     515] = 32'h78a62e2a;
    ram_cell[     516] = 32'h0d659beb;
    ram_cell[     517] = 32'hd7b94690;
    ram_cell[     518] = 32'hf5c0481b;
    ram_cell[     519] = 32'h183ced36;
    ram_cell[     520] = 32'haf31400a;
    ram_cell[     521] = 32'hf2a8c6d2;
    ram_cell[     522] = 32'hec9ce9b8;
    ram_cell[     523] = 32'h40a63fa2;
    ram_cell[     524] = 32'h3626007b;
    ram_cell[     525] = 32'hf67d9176;
    ram_cell[     526] = 32'h0a4b4fdc;
    ram_cell[     527] = 32'ha72dbd86;
    ram_cell[     528] = 32'h62c3d056;
    ram_cell[     529] = 32'hc301581a;
    ram_cell[     530] = 32'h392c32c0;
    ram_cell[     531] = 32'hf9092a1b;
    ram_cell[     532] = 32'haed2e2fe;
    ram_cell[     533] = 32'hfa29828c;
    ram_cell[     534] = 32'hf92c4a12;
    ram_cell[     535] = 32'he55a5672;
    ram_cell[     536] = 32'h00edd8b3;
    ram_cell[     537] = 32'hbdbaeaf9;
    ram_cell[     538] = 32'h08d3b198;
    ram_cell[     539] = 32'h200de9ee;
    ram_cell[     540] = 32'h7e6f3ae0;
    ram_cell[     541] = 32'hee865c7e;
    ram_cell[     542] = 32'h6dae476c;
    ram_cell[     543] = 32'haa37a9a7;
    ram_cell[     544] = 32'hea17086c;
    ram_cell[     545] = 32'hf4b074b2;
    ram_cell[     546] = 32'h67145e39;
    ram_cell[     547] = 32'hee54e980;
    ram_cell[     548] = 32'h09114575;
    ram_cell[     549] = 32'h6d6160a7;
    ram_cell[     550] = 32'hd986764a;
    ram_cell[     551] = 32'h19543bff;
    ram_cell[     552] = 32'he529bad1;
    ram_cell[     553] = 32'hdb905c3a;
    ram_cell[     554] = 32'hee654517;
    ram_cell[     555] = 32'h6e7ba4a1;
    ram_cell[     556] = 32'h7ded65a3;
    ram_cell[     557] = 32'hd79bc35c;
    ram_cell[     558] = 32'h9cfaddc3;
    ram_cell[     559] = 32'h89c74c71;
    ram_cell[     560] = 32'h4c76a75f;
    ram_cell[     561] = 32'h61d3cf3c;
    ram_cell[     562] = 32'hff770b0c;
    ram_cell[     563] = 32'he1825087;
    ram_cell[     564] = 32'hdfa74abd;
    ram_cell[     565] = 32'hc16e441c;
    ram_cell[     566] = 32'h69047953;
    ram_cell[     567] = 32'h5f410200;
    ram_cell[     568] = 32'h9dec90e6;
    ram_cell[     569] = 32'h18ae62c9;
    ram_cell[     570] = 32'h4ffbfbfb;
    ram_cell[     571] = 32'h7a7f0d72;
    ram_cell[     572] = 32'h48448d0d;
    ram_cell[     573] = 32'hcd4791a8;
    ram_cell[     574] = 32'h5a72ad43;
    ram_cell[     575] = 32'hd7ed9c6d;
    ram_cell[     576] = 32'h91942cb9;
    ram_cell[     577] = 32'h43a6496d;
    ram_cell[     578] = 32'he580c72c;
    ram_cell[     579] = 32'h311b363f;
    ram_cell[     580] = 32'h87907a90;
    ram_cell[     581] = 32'h2b21a413;
    ram_cell[     582] = 32'h53b8e1d6;
    ram_cell[     583] = 32'h88250a32;
    ram_cell[     584] = 32'h09c5a37a;
    ram_cell[     585] = 32'hc2243a91;
    ram_cell[     586] = 32'ha1693490;
    ram_cell[     587] = 32'h191748dc;
    ram_cell[     588] = 32'h2992ae1f;
    ram_cell[     589] = 32'hc63d4890;
    ram_cell[     590] = 32'h8ccecd70;
    ram_cell[     591] = 32'h3193708d;
    ram_cell[     592] = 32'h913e3775;
    ram_cell[     593] = 32'hd910e426;
    ram_cell[     594] = 32'hcc26feb9;
    ram_cell[     595] = 32'heb0eeeba;
    ram_cell[     596] = 32'h9a50a17b;
    ram_cell[     597] = 32'h80b84775;
    ram_cell[     598] = 32'h3f97149d;
    ram_cell[     599] = 32'hf6ac474b;
    ram_cell[     600] = 32'h992a07b3;
    ram_cell[     601] = 32'h445da2b4;
    ram_cell[     602] = 32'hafe7eb6a;
    ram_cell[     603] = 32'h90bceed3;
    ram_cell[     604] = 32'h71359bc6;
    ram_cell[     605] = 32'h128c3e13;
    ram_cell[     606] = 32'h78d55076;
    ram_cell[     607] = 32'h7aadd851;
    ram_cell[     608] = 32'hd5b022ae;
    ram_cell[     609] = 32'h4964f1b4;
    ram_cell[     610] = 32'hc375138b;
    ram_cell[     611] = 32'hb85e82c8;
    ram_cell[     612] = 32'h218ba89d;
    ram_cell[     613] = 32'ha70b2663;
    ram_cell[     614] = 32'haeb1df6c;
    ram_cell[     615] = 32'h44c72fc9;
    ram_cell[     616] = 32'he6a6c5bc;
    ram_cell[     617] = 32'h6cfb186d;
    ram_cell[     618] = 32'h22891f8d;
    ram_cell[     619] = 32'h0a6d0ae0;
    ram_cell[     620] = 32'h9b14b6bb;
    ram_cell[     621] = 32'h5f9787a9;
    ram_cell[     622] = 32'hf5abf036;
    ram_cell[     623] = 32'h8cfad753;
    ram_cell[     624] = 32'hdf4bfef5;
    ram_cell[     625] = 32'h3d35a948;
    ram_cell[     626] = 32'hb9bc0ce9;
    ram_cell[     627] = 32'h57a77477;
    ram_cell[     628] = 32'h70dce3d0;
    ram_cell[     629] = 32'he4e2830f;
    ram_cell[     630] = 32'h8c620401;
    ram_cell[     631] = 32'hef713af2;
    ram_cell[     632] = 32'h14d0ce4c;
    ram_cell[     633] = 32'h109ef8cf;
    ram_cell[     634] = 32'h4138cfbb;
    ram_cell[     635] = 32'h87e88988;
    ram_cell[     636] = 32'h61bbf763;
    ram_cell[     637] = 32'hf9fa2463;
    ram_cell[     638] = 32'ha7f8399d;
    ram_cell[     639] = 32'hb142b2b5;
    ram_cell[     640] = 32'h865839cc;
    ram_cell[     641] = 32'h61b25842;
    ram_cell[     642] = 32'h80d22ca5;
    ram_cell[     643] = 32'h0f9b2848;
    ram_cell[     644] = 32'hf8230e0d;
    ram_cell[     645] = 32'h18a3b981;
    ram_cell[     646] = 32'h9eb016a3;
    ram_cell[     647] = 32'h059b7f34;
    ram_cell[     648] = 32'h9e13f060;
    ram_cell[     649] = 32'h4d285998;
    ram_cell[     650] = 32'h712a4809;
    ram_cell[     651] = 32'heea4d035;
    ram_cell[     652] = 32'h81463bcd;
    ram_cell[     653] = 32'h25612af6;
    ram_cell[     654] = 32'ha915f294;
    ram_cell[     655] = 32'h9a8b3f89;
    ram_cell[     656] = 32'h4a9bfe3b;
    ram_cell[     657] = 32'h3f1032d1;
    ram_cell[     658] = 32'h740f6701;
    ram_cell[     659] = 32'h76d6e490;
    ram_cell[     660] = 32'h67aee858;
    ram_cell[     661] = 32'hca0e8ba5;
    ram_cell[     662] = 32'h0c47e961;
    ram_cell[     663] = 32'hfdf4aac8;
    ram_cell[     664] = 32'hec81780c;
    ram_cell[     665] = 32'h7db13aad;
    ram_cell[     666] = 32'hc9e20e69;
    ram_cell[     667] = 32'h8b61c48b;
    ram_cell[     668] = 32'hc16c8a42;
    ram_cell[     669] = 32'hd9c61fa7;
    ram_cell[     670] = 32'he1d594bd;
    ram_cell[     671] = 32'h3c6ad86e;
    ram_cell[     672] = 32'h9f102443;
    ram_cell[     673] = 32'h9307829d;
    ram_cell[     674] = 32'hd34dfc84;
    ram_cell[     675] = 32'h00f27d40;
    ram_cell[     676] = 32'h9bf68f08;
    ram_cell[     677] = 32'hbf22ac6a;
    ram_cell[     678] = 32'hf1c8acdf;
    ram_cell[     679] = 32'h5df3549e;
    ram_cell[     680] = 32'h0e3759a5;
    ram_cell[     681] = 32'h75a18a3e;
    ram_cell[     682] = 32'hed3e8f54;
    ram_cell[     683] = 32'hb8dfe335;
    ram_cell[     684] = 32'h00a00725;
    ram_cell[     685] = 32'hd75c57d4;
    ram_cell[     686] = 32'hf42e0ccd;
    ram_cell[     687] = 32'hf91930d7;
    ram_cell[     688] = 32'hb7cb9e13;
    ram_cell[     689] = 32'h1cc57d47;
    ram_cell[     690] = 32'hc31c72e6;
    ram_cell[     691] = 32'h3f56ec06;
    ram_cell[     692] = 32'h61f9446d;
    ram_cell[     693] = 32'h7627294f;
    ram_cell[     694] = 32'h5652bf23;
    ram_cell[     695] = 32'h046aac35;
    ram_cell[     696] = 32'h105222d7;
    ram_cell[     697] = 32'he6b1f975;
    ram_cell[     698] = 32'h8ca9a1a6;
    ram_cell[     699] = 32'h1b8731be;
    ram_cell[     700] = 32'h2768821c;
    ram_cell[     701] = 32'h7248a000;
    ram_cell[     702] = 32'he39b99a5;
    ram_cell[     703] = 32'h5ea64d5c;
    ram_cell[     704] = 32'h81bd980b;
    ram_cell[     705] = 32'hd7937f6e;
    ram_cell[     706] = 32'h3a879af8;
    ram_cell[     707] = 32'h38e3e264;
    ram_cell[     708] = 32'h3b14c1a1;
    ram_cell[     709] = 32'hacc93abd;
    ram_cell[     710] = 32'h00633e22;
    ram_cell[     711] = 32'h2af068d5;
    ram_cell[     712] = 32'h0243964a;
    ram_cell[     713] = 32'hc00bd7eb;
    ram_cell[     714] = 32'hf00d50e5;
    ram_cell[     715] = 32'h9bba1f72;
    ram_cell[     716] = 32'h6a3160e2;
    ram_cell[     717] = 32'hf3c15358;
    ram_cell[     718] = 32'h11fae70b;
    ram_cell[     719] = 32'h766bd2b9;
    ram_cell[     720] = 32'hab683272;
    ram_cell[     721] = 32'h4d2cf791;
    ram_cell[     722] = 32'h1821e334;
    ram_cell[     723] = 32'h6dc93f79;
    ram_cell[     724] = 32'h0bc22f81;
    ram_cell[     725] = 32'h32064f41;
    ram_cell[     726] = 32'h01c8d4d5;
    ram_cell[     727] = 32'h0e220c87;
    ram_cell[     728] = 32'h369ae6a8;
    ram_cell[     729] = 32'h8ce1cb93;
    ram_cell[     730] = 32'h7777a300;
    ram_cell[     731] = 32'h15634e56;
    ram_cell[     732] = 32'hefdb8f44;
    ram_cell[     733] = 32'h2f209ac4;
    ram_cell[     734] = 32'heea97b8c;
    ram_cell[     735] = 32'h3ddc1664;
    ram_cell[     736] = 32'h6a120c94;
    ram_cell[     737] = 32'h7e9eb747;
    ram_cell[     738] = 32'hb36909b1;
    ram_cell[     739] = 32'h49c8d695;
    ram_cell[     740] = 32'h652c0f39;
    ram_cell[     741] = 32'hf0ad54c8;
    ram_cell[     742] = 32'he27cc0d1;
    ram_cell[     743] = 32'h7ad81008;
    ram_cell[     744] = 32'h5aa3b537;
    ram_cell[     745] = 32'hc634a896;
    ram_cell[     746] = 32'hbfb98720;
    ram_cell[     747] = 32'h6fdd74be;
    ram_cell[     748] = 32'hf4de52c3;
    ram_cell[     749] = 32'hf51565ff;
    ram_cell[     750] = 32'h628ec3a8;
    ram_cell[     751] = 32'hc3d211e6;
    ram_cell[     752] = 32'h1020e580;
    ram_cell[     753] = 32'hea85bdb3;
    ram_cell[     754] = 32'h58c16785;
    ram_cell[     755] = 32'h20424dc4;
    ram_cell[     756] = 32'h17764283;
    ram_cell[     757] = 32'h328a996b;
    ram_cell[     758] = 32'h16c4a699;
    ram_cell[     759] = 32'hbddcf060;
    ram_cell[     760] = 32'h7c2c3516;
    ram_cell[     761] = 32'h87538398;
    ram_cell[     762] = 32'h3cf4bdf7;
    ram_cell[     763] = 32'hd506e2bf;
    ram_cell[     764] = 32'hc4fcb614;
    ram_cell[     765] = 32'hb381e0f2;
    ram_cell[     766] = 32'hb52483a5;
    ram_cell[     767] = 32'hf46409c2;
end

endmodule

